magic
tech sky130A
timestamp 1719085816
<< metal1 >>
rect 326 -1365 362 -1361
rect 326 -1453 330 -1365
rect 357 -1453 362 -1365
rect 326 -1457 362 -1453
<< via1 >>
rect 330 -1453 357 -1365
<< metal2 >>
rect 326 -1365 362 -1361
rect 326 -1453 330 -1365
rect 357 -1453 362 -1365
rect 326 -1457 362 -1453
<< end >>
