magic
tech sky130A
magscale 1 2
timestamp 1719091984
<< dnwell >>
rect 683 -653 5288 1461
rect 683 -659 2069 -653
<< nwell >>
rect 573 1255 5397 1570
rect 573 -447 769 1255
rect 5082 -447 5397 1255
rect 573 -762 5397 -447
<< mvnsubdiff >>
rect 640 1484 5331 1504
rect 640 1450 720 1484
rect 5251 1450 5331 1484
rect 640 1430 5331 1450
rect 640 1424 714 1430
rect 640 -616 660 1424
rect 694 -616 714 1424
rect 640 -622 714 -616
rect 5257 1424 5331 1430
rect 5257 -616 5277 1424
rect 5311 -616 5331 1424
rect 5257 -622 5331 -616
rect 640 -642 5331 -622
rect 640 -676 720 -642
rect 5251 -676 5331 -642
rect 640 -696 5331 -676
<< mvnsubdiffcont >>
rect 720 1450 5251 1484
rect 660 -616 694 1424
rect 5277 -616 5311 1424
rect 720 -676 5251 -642
<< locali >>
rect 660 1450 720 1484
rect 5251 1450 5311 1484
rect 660 1424 5311 1450
rect 694 1348 5277 1424
rect 694 1305 881 1348
rect 694 -246 777 1305
rect 820 1263 881 1305
rect 3560 1276 5028 1286
rect 820 1255 2950 1263
rect 820 1220 1062 1255
rect 2925 1220 2950 1255
rect 820 1169 2950 1220
rect 3560 1230 3582 1276
rect 5010 1230 5028 1276
rect 3560 1196 5028 1230
rect 820 465 881 1169
rect 4868 1166 4994 1196
rect 820 436 2960 465
rect 4868 458 4914 1166
rect 820 373 871 436
rect 2899 373 2960 436
rect 820 345 2960 373
rect 3679 436 4914 458
rect 3679 379 3742 436
rect 4827 379 4914 436
rect 3679 351 4914 379
rect 820 -246 881 345
rect 694 -353 881 -246
rect 4868 -331 4914 351
rect 4970 -331 4994 1166
rect 4868 -345 4994 -331
rect 694 -374 2963 -353
rect 694 -431 903 -374
rect 2929 -431 2963 -374
rect 694 -453 2963 -431
rect 3560 -407 5063 -345
rect 3560 -444 3603 -407
rect 5003 -444 5063 -407
rect 694 -542 881 -453
rect 3560 -462 5063 -444
rect 5126 -542 5277 1348
rect 694 -616 5277 -542
rect 660 -642 5311 -616
rect 660 -676 720 -642
rect 5251 -676 5311 -642
<< viali >>
rect 777 -246 820 1305
rect 1062 1220 2925 1255
rect 3582 1230 5010 1276
rect 871 373 2899 436
rect 3742 379 4827 436
rect 4914 -331 4970 1166
rect 903 -431 2929 -374
rect 3603 -444 5003 -407
<< metal1 >>
rect 3194 1386 3262 1567
rect 3334 1386 3402 1567
rect 3475 1390 3542 1566
rect 761 1332 881 1333
rect 761 1308 3152 1332
rect 761 1305 1088 1308
rect 761 -246 777 1305
rect 820 1255 1088 1305
rect 820 1220 1062 1255
rect 820 1194 1088 1220
rect 2943 1194 3152 1308
rect 820 1186 3152 1194
rect 820 465 881 1186
rect 3208 1092 3248 1386
rect 1023 1046 3248 1092
rect 3003 564 3049 1046
rect 3348 960 3384 1386
rect 3486 1075 3522 1390
rect 3554 1276 5081 1332
rect 3554 1230 3582 1276
rect 5010 1230 5081 1276
rect 3554 1186 5081 1230
rect 4868 1166 4994 1186
rect 3486 1030 4784 1075
rect 3602 1029 4784 1030
rect 3602 1000 3649 1029
rect 3348 924 3474 960
rect 3438 574 3474 924
rect 1027 518 3049 564
rect 820 436 2960 465
rect 820 373 871 436
rect 2899 373 2960 436
rect 820 345 2960 373
rect 820 -246 881 345
rect 3003 291 3049 518
rect 1027 245 3049 291
rect 3003 -237 3049 245
rect 761 -356 881 -246
rect 1031 -265 3049 -237
rect 3179 512 3287 517
rect 3179 501 3362 512
rect 3179 327 3188 501
rect 3278 327 3362 501
rect 3179 312 3362 327
rect 1031 -283 3047 -265
rect 3179 -356 3287 312
rect 3442 256 3470 574
rect 3601 568 3649 1000
rect 3601 519 4780 568
rect 3601 289 3649 519
rect 4868 458 4914 1166
rect 3679 436 4914 458
rect 3679 379 3742 436
rect 4827 379 4914 436
rect 3679 351 4914 379
rect 3601 243 4784 289
rect 3601 -221 3649 243
rect 3601 -266 4784 -221
rect 3603 -267 4784 -266
rect 4868 -331 4914 351
rect 4970 -331 4994 1166
rect 4868 -356 4994 -331
rect 761 -374 3062 -356
rect 761 -431 903 -374
rect 2929 -431 3062 -374
rect 761 -502 3062 -431
rect 3179 -380 5063 -356
rect 3179 -495 3419 -380
rect 5008 -495 5063 -380
rect 3179 -502 5063 -495
<< via1 >>
rect 1088 1255 2943 1308
rect 1088 1220 2925 1255
rect 2925 1220 2943 1255
rect 1088 1194 2943 1220
rect 3188 327 3278 501
rect 3419 -407 5008 -380
rect 3419 -444 3603 -407
rect 3603 -444 5003 -407
rect 5003 -444 5008 -407
rect 3419 -495 5008 -444
<< metal2 >>
rect 735 1308 5169 1336
rect 735 1194 1088 1308
rect 2943 1194 5169 1308
rect 735 1141 5169 1194
rect 4886 1016 5062 1023
rect 961 824 5062 1016
rect 4886 823 5062 824
rect 961 584 4813 776
rect 3179 501 3360 509
rect 3179 327 3188 501
rect 3278 327 3360 501
rect 3179 319 3360 327
rect 3450 235 3647 584
rect 961 43 4813 235
rect 4886 -17 5062 -9
rect 961 -209 5062 -17
rect 726 -380 5160 -331
rect 726 -495 3419 -380
rect 5008 -495 5160 -380
rect 726 -526 5160 -495
use iso_switch_via  iso_switch_via_0
timestamp 1719085816
transform 1 0 3912 0 1 2722
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_1
timestamp 1719085816
transform 1 0 625 0 1 2709
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_2
timestamp 1719085816
transform 1 0 1100 0 1 2938
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_3
timestamp 1719085816
transform 1 0 1257 0 1 2709
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_4
timestamp 1719085816
transform 1 0 1573 0 1 2709
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_5
timestamp 1719085816
transform 1 0 1889 0 1 2709
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_6
timestamp 1719085816
transform 1 0 945 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_7
timestamp 1719085816
transform 1 0 2205 0 1 2709
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_8
timestamp 1719085816
transform 1 0 468 0 1 2938
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_9
timestamp 1719085816
transform 1 0 784 0 1 2938
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_10
timestamp 1719085816
transform 1 0 2048 0 1 2938
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_11
timestamp 1719085816
transform 1 0 1416 0 1 2938
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_12
timestamp 1719085816
transform 1 0 1732 0 1 2938
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_13
timestamp 1719085816
transform 1 0 629 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_14
timestamp 1719085816
transform 1 0 1100 0 -1 -1898
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_15
timestamp 1719085816
transform 1 0 1261 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_16
timestamp 1719085816
transform 1 0 1577 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_17
timestamp 1719085816
transform 1 0 309 0 1 2705
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_18
timestamp 1719085816
transform 1 0 1893 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_19
timestamp 1719085816
transform 1 0 2209 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_20
timestamp 1719085816
transform 1 0 941 0 1 2709
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_21
timestamp 1719085816
transform 1 0 468 0 -1 -1898
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_22
timestamp 1719085816
transform 1 0 784 0 -1 -1898
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_23
timestamp 1719085816
transform 1 0 2048 0 -1 -1898
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_24
timestamp 1719085816
transform 1 0 1416 0 -1 -1898
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_25
timestamp 1719085816
transform 1 0 1732 0 -1 -1898
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_26
timestamp 1719085816
transform 1 0 3280 0 1 2722
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_27
timestamp 1719085816
transform -1 0 4494 0 1 2934
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_28
timestamp 1719085816
transform 1 0 3596 0 1 2722
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_29
timestamp 1719085816
transform -1 0 4810 0 1 2934
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_30
timestamp 1719085816
transform -1 0 5126 0 1 2934
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_31
timestamp 1719085816
transform -1 0 5442 0 1 3722
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_32
timestamp 1719085816
transform 1 0 3912 0 1 3510
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_33
timestamp 1719085816
transform -1 0 5126 0 1 3722
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_34
timestamp 1719085816
transform -1 0 5442 0 1 2934
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_35
timestamp 1719085816
transform 1 0 3596 0 1 3510
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_36
timestamp 1719085816
transform -1 0 4054 0 1 3234
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_37
timestamp 1719085816
transform -1 0 4222 0 1 3235
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_38
timestamp 1719085816
transform 1 0 309 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_39
timestamp 1719085816
transform -1 0 4810 0 1 3722
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_40
timestamp 1719085816
transform 1 0 3280 0 1 3510
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_41
timestamp 1719085816
transform -1 0 4494 0 1 3722
box 652 -2914 724 -2722
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  sky130_fd_pr__nfet_g5v0d10v5_EJGQJV_0 paramcells
timestamp 1719085816
transform -1 0 3456 0 1 412
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_SABQJA  sky130_fd_pr__nfet_g5v0d10v5_SABQJA_0 paramcells
timestamp 1719083619
transform -1 0 4282 0 1 11
box -673 -458 673 458
use sky130_fd_pr__pfet_g5v0d10v5_LQS9ZD  sky130_fd_pr__pfet_g5v0d10v5_LQS9ZD_0 paramcells
timestamp 1719083619
transform 1 0 1946 0 1 4
box -1177 -497 1177 497
use sky130_fd_pr__pfet_g5v0d10v5_LQS9ZD  XM4
timestamp 1719083619
transform 1 0 1946 0 1 808
box -1177 -497 1177 497
use sky130_fd_pr__nfet_g5v0d10v5_SABQJA  XM15
timestamp 1719083619
transform -1 0 4282 0 1 797
box -673 -458 673 458
<< labels >>
flabel metal2 4886 -209 5062 -9 0 FreeSans 256 180 0 0 out
port 3 nsew
flabel metal2 4886 823 5062 1023 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal1 3334 1386 3402 1567 0 FreeSans 256 270 0 0 shunt
port 6 nsew
flabel metal1 845 1186 1045 1264 0 FreeSans 256 0 0 0 vdd
port 5 nsew
flabel metal1 3475 1390 3542 1566 0 FreeSans 256 270 0 0 on
port 0 nsew
flabel metal1 3194 1386 3262 1567 0 FreeSans 256 270 0 0 off
port 1 nsew
flabel metal1 3180 -463 3380 -356 0 FreeSans 256 180 0 0 vss
port 2 nsew
<< end >>
