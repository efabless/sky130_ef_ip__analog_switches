** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch_ena1v8.sch
.subckt simple_analog_switch_ena1v8 avss on out in avdd dvdd dvss
*.PININFO on:I avss:B out:B in:B avdd:B dvdd:B dvss:B
x2 on dvdd dvss dvss avdd avdd net3 sky130_fd_sc_hvl__lsbuflv2hv_1
XD1 dvss on sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
x3 net1 net2 avss out in avdd simple_analog_switch
x1 net3 dvss dvss avdd avdd net2 sky130_fd_sc_hvl__inv_2
x4 net2 dvss dvss avdd avdd net1 sky130_fd_sc_hvl__inv_2
x5[1] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
x5[0] dvss dvss avdd avdd sky130_fd_sc_hvl__decap_4
.ends

* expanding   symbol:  simple_analog_switch.sym # of pins=6
** sym_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch.sym
** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_ef_ip__analog_switches/xschem/simple_analog_switch.sch
.subckt simple_analog_switch on off vss out in vdd
*.PININFO on:I out:B vdd:B vss:B in:B off:I
XM1 in on out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
XM2 in off out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=8 nf=4 m=1
XM3 out off out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM4 out on out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
XM5 in off in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM6 in on in vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
.ends

.end
