magic
tech sky130A
magscale 1 2
timestamp 1716605065
<< psubdiff >>
rect 41 1640 65 1724
rect 4354 1640 4378 1724
<< psubdiffcont >>
rect 65 1640 4354 1724
<< locali >>
rect 2566 3229 2629 3295
rect 2879 3275 3095 3283
rect 2879 3230 2890 3275
rect 3085 3230 3095 3275
rect 2879 3221 3095 3230
rect 756 2379 996 2392
rect 756 2337 770 2379
rect 982 2337 996 2379
rect 756 2324 996 2337
rect 2444 2347 2684 2353
rect 2444 2295 2460 2347
rect 2668 2295 2684 2347
rect 2444 2287 2684 2295
rect 2851 2348 3091 2354
rect 2851 2296 2867 2348
rect 3075 2296 3091 2348
rect 2851 2288 3091 2296
rect 352 2048 408 2056
rect 352 1964 360 2048
rect 398 1994 408 2048
rect 398 1964 492 1994
rect 352 1960 492 1964
rect 352 1954 408 1960
rect 49 1640 65 1724
rect 4354 1640 4370 1724
<< viali >>
rect 2890 3230 3085 3275
rect 770 2337 982 2379
rect 2460 2295 2668 2347
rect 2867 2296 3075 2348
rect 360 1964 398 2048
rect 1009 1640 1199 1724
<< metal1 >>
rect 0 3604 498 3627
rect 1001 3619 1208 3628
rect 1001 3604 1011 3619
rect 0 3538 1011 3604
rect 0 3479 498 3538
rect 1001 3490 1011 3538
rect 1198 3604 1208 3619
rect 1198 3538 3461 3604
rect 1198 3490 1208 3538
rect 1001 3480 1208 3490
rect 2869 3275 3111 3283
rect 2869 3230 2890 3275
rect 3085 3230 3111 3275
rect 2869 3221 3111 3230
rect 615 2903 837 2916
rect 615 2868 627 2903
rect 491 2730 627 2868
rect 615 2677 627 2730
rect 826 2868 837 2903
rect 1804 2903 2027 2916
rect 1804 2868 1816 2903
rect 826 2730 1816 2868
rect 826 2677 837 2730
rect 615 2666 837 2677
rect 1804 2678 1816 2730
rect 2013 2868 2027 2903
rect 2013 2730 3464 2868
rect 2013 2678 2027 2730
rect 1804 2666 2027 2678
rect 1 2581 517 2638
rect 1 2530 263 2581
rect 756 2379 996 2392
rect 756 2365 770 2379
rect 403 2337 770 2365
rect 982 2337 996 2379
rect 403 2329 996 2337
rect 2 2129 289 2130
rect 403 2129 439 2329
rect 756 2324 996 2329
rect 2444 2347 2684 2353
rect 2444 2295 2460 2347
rect 2668 2295 2684 2347
rect 2444 2287 2684 2295
rect 2851 2348 3091 2354
rect 2851 2296 2867 2348
rect 3075 2296 3091 2348
rect 2851 2288 3091 2296
rect 2 2093 439 2129
rect 2 2041 289 2093
rect 348 2048 3468 2056
rect 348 1964 360 2048
rect 398 1980 3468 2048
rect 398 1964 496 1980
rect 348 1954 496 1964
rect 996 1724 1213 1735
rect 996 1640 1009 1724
rect 1199 1640 1213 1724
rect 996 1630 1213 1640
rect 0 1162 273 1308
rect 615 1302 837 1308
rect 615 1169 624 1302
rect 830 1169 837 1302
rect 615 1162 837 1169
rect 1805 1301 2027 1308
rect 1805 1170 1814 1301
rect 2019 1170 2027 1301
rect 1805 1162 2027 1170
rect 0 260 255 406
<< via1 >>
rect 1011 3490 1198 3619
rect 627 2677 826 2903
rect 1816 2678 2013 2903
rect 1009 1640 1199 1724
rect 624 1169 830 1302
rect 1814 1170 2019 1301
<< metal2 >>
rect 1001 3619 1208 3628
rect 1001 3490 1011 3619
rect 1198 3490 1208 3619
rect 615 2903 837 2916
rect 615 2677 627 2903
rect 826 2677 837 2903
rect 615 1302 837 2677
rect 1001 1724 1208 3490
rect 1804 2903 2027 2916
rect 1804 2678 1816 2903
rect 2013 2678 2027 2903
rect 2883 2813 2931 3252
rect 1804 2666 2027 2678
rect 1001 1640 1009 1724
rect 1199 1640 1208 1724
rect 1001 1630 1208 1640
rect 615 1169 624 1302
rect 830 1169 837 1302
rect 615 1162 837 1169
rect 1805 1301 2027 2666
rect 2626 2765 2931 2813
rect 2626 2491 2674 2765
rect 2626 2443 3206 2491
rect 2626 2283 2674 2443
rect 2816 2358 2883 2359
rect 2801 2287 2883 2358
rect 2958 2287 3006 2295
rect 2801 2202 2851 2287
rect 2418 2152 2851 2202
rect 2418 1540 2468 2152
rect 3158 2024 3206 2443
rect 2523 1976 3206 2024
rect 2523 1526 2571 1976
rect 1805 1170 1814 1301
rect 2019 1170 2027 1301
rect 1805 1162 2027 1170
rect 4118 800 4416 1000
rect 4119 561 4416 760
use iso_switch_via  iso_switch_via_0
timestamp 1716604942
transform 0 1 5797 1 0 2564
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_1
timestamp 1716604942
transform 0 1 5380 1 0 1630
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_2
timestamp 1716604942
transform 0 1 5797 1 0 1635
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_3
timestamp 1716604942
transform -1 0 3130 0 1 4282
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_13
timestamp 1716604942
transform -1 0 3235 0 1 4277
box 652 -2914 724 -2722
use simple_analog_switch  simple_analog_switch_0
timestamp 1716604942
transform 1 0 -577 0 1 -24
box 577 24 4993 1570
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  sky130_fd_pr__diode_pw2nd_05v5_FT76RJ_0 paramcells
timestamp 1716604942
transform 1 0 239 0 1 2082
box -183 -183 183 183
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1716604942
transform 1 0 3083 0 -1 3605
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_1
timestamp 1716604942
transform 1 0 3083 0 1 1977
box -66 -43 450 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1716604942
transform 1 0 2603 0 1 1977
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_1
timestamp 1716604942
transform 1 0 2603 0 -1 3605
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1716604942
transform 1 0 491 0 1 1977
box -66 -43 2178 1671
<< labels >>
flabel locali s 3041 2294 3075 2328 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel metal1 0 1162 156 1308 0 FreeSans 800 0 0 0 avdd
port 4 nsew
flabel metal1 0 260 156 406 0 FreeSans 800 0 0 0 avss
port 5 nsew
flabel metal1 1 2530 263 2638 0 FreeSans 800 0 0 0 dvdd
port 6 nsew
flabel metal1 0 3479 263 3627 0 FreeSans 800 0 0 0 dvss
port 7 nsew
flabel metal1 2 2041 182 2130 0 FreeSans 800 0 0 0 on
port 8 nsew
flabel metal2 4230 800 4416 1000 0 FreeSans 800 0 0 0 in
port 2 nsew
flabel metal2 4230 561 4416 760 0 FreeSans 800 0 0 0 out
port 3 nsew
<< end >>
