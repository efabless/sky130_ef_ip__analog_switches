magic
tech sky130A
magscale 1 2
timestamp 1724439637
<< psubdiff >>
rect 61 1640 85 1724
rect 3514 1640 3538 1724
<< psubdiffcont >>
rect 85 1640 3514 1724
<< locali >>
rect 2566 3229 2629 3295
rect 2879 3275 3095 3283
rect 2879 3230 2890 3275
rect 3085 3230 3095 3275
rect 2879 3221 3095 3230
rect 756 2379 996 2392
rect 756 2337 770 2379
rect 982 2337 996 2379
rect 756 2324 996 2337
rect 2444 2347 2684 2353
rect 2444 2295 2460 2347
rect 2668 2295 2684 2347
rect 2444 2287 2684 2295
rect 2851 2348 3091 2354
rect 2851 2296 2867 2348
rect 3075 2296 3091 2348
rect 2851 2288 3091 2296
rect 69 1640 85 1724
rect 3514 1640 3530 1724
rect 612 1454 844 1466
rect 612 1414 624 1454
rect 830 1414 844 1454
rect 612 1400 844 1414
<< viali >>
rect 2890 3230 3085 3275
rect 770 2337 982 2379
rect 380 2147 426 2302
rect 2460 2295 2668 2347
rect 2867 2296 3075 2348
rect 1009 1640 1199 1724
rect 624 1414 830 1454
<< metal1 >>
rect 0 3604 498 3627
rect 0 3559 3461 3604
rect 0 3538 1011 3559
rect 0 3479 498 3538
rect 1001 3430 1011 3538
rect 1198 3538 3461 3559
rect 1198 3430 1208 3538
rect 1001 3420 1208 3430
rect 2869 3275 3111 3283
rect 2869 3230 2890 3275
rect 3085 3230 3111 3275
rect 2869 3221 3111 3230
rect 615 2903 837 2916
rect 615 2868 627 2903
rect 299 2730 627 2868
rect 615 2677 627 2730
rect 826 2868 837 2903
rect 1543 2903 1766 2916
rect 1543 2868 1555 2903
rect 826 2730 1555 2868
rect 826 2677 837 2730
rect 615 2666 837 2677
rect 1543 2678 1555 2730
rect 1752 2868 1766 2903
rect 1752 2730 3464 2868
rect 1752 2678 1766 2730
rect 1543 2666 1766 2678
rect 1 2581 517 2638
rect 1 2530 263 2581
rect 756 2379 996 2392
rect 756 2365 770 2379
rect 367 2337 770 2365
rect 982 2337 996 2379
rect 367 2329 996 2337
rect 367 2302 439 2329
rect 756 2324 996 2329
rect 2444 2347 2684 2353
rect 367 2169 380 2302
rect 223 2147 380 2169
rect 426 2147 439 2302
rect 2444 2295 2460 2347
rect 2668 2295 2684 2347
rect 2444 2287 2684 2295
rect 2851 2348 3091 2354
rect 2851 2296 2867 2348
rect 3075 2296 3091 2348
rect 2851 2288 3091 2296
rect 223 2133 439 2147
rect 223 2130 262 2133
rect 2 2041 262 2130
rect 299 1980 1010 2056
rect 1200 1980 3468 2056
rect 996 1724 1213 1735
rect 996 1640 1009 1724
rect 1199 1640 1213 1724
rect 996 1630 1213 1640
rect 612 1464 844 1466
rect 612 1410 624 1464
rect 832 1410 844 1464
rect 612 1400 844 1410
rect 604 1302 1804 1310
rect 604 1169 624 1302
rect 1795 1169 1804 1302
rect 604 1166 1804 1169
rect 615 1162 837 1166
<< via1 >>
rect 1011 3430 1198 3559
rect 627 2677 826 2903
rect 1555 2678 1752 2903
rect 1010 1968 1200 2094
rect 1009 1640 1199 1724
rect 624 1454 832 1464
rect 624 1414 830 1454
rect 830 1414 832 1454
rect 624 1410 832 1414
rect 624 1169 1795 1302
rect 2060 -322 3191 -198
<< metal2 >>
rect 1001 3559 1208 3568
rect 1001 3430 1011 3559
rect 1198 3430 1208 3559
rect 615 2903 837 2916
rect 615 2677 627 2903
rect 826 2677 837 2903
rect 615 1464 837 2677
rect 1001 2094 1208 3430
rect 1001 1968 1010 2094
rect 1200 1968 1208 2094
rect 1001 1724 1208 1968
rect 1001 1640 1009 1724
rect 1199 1640 1208 1724
rect 1001 1630 1208 1640
rect 1543 2903 1766 2916
rect 1543 2678 1555 2903
rect 1752 2678 1766 2903
rect 2883 2813 2931 3252
rect 1543 2658 1766 2678
rect 2626 2765 2931 2813
rect 615 1410 624 1464
rect 832 1410 837 1464
rect 615 1310 837 1410
rect 1543 1310 1765 2658
rect 1845 2304 2487 2354
rect 1845 1540 1895 2304
rect 2626 2283 2674 2765
rect 2816 2358 2883 2359
rect 2801 2287 2883 2358
rect 2958 2287 3006 2295
rect 2801 2202 2851 2287
rect 1950 2152 2851 2202
rect 1950 1526 1998 2152
rect -4 1302 3500 1310
rect -4 1169 624 1302
rect 1795 1169 3500 1302
rect -4 1120 3500 1169
rect 3196 540 3494 972
rect 3197 -20 3495 412
rect 0 -198 3482 -172
rect 0 -322 2060 -198
rect 3191 -322 3482 -198
rect 0 -340 3482 -322
use iso_switch_via  iso_switch_via_0
timestamp 1719085816
transform 0 1 5797 1 0 2564
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_1
timestamp 1719085816
transform 0 1 5380 1 0 1630
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_2
timestamp 1719085816
transform 0 1 5797 1 0 1635
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_3
timestamp 1719085816
transform -1 0 2557 0 1 4282
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_13
timestamp 1719085816
transform -1 0 2662 0 1 4277
box 652 -2914 724 -2722
use simple_analog_switch_2  simple_analog_switch_2_0
timestamp 1724439637
transform 1 0 -1149 0 1 -624
box 1210 24 4680 2170
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1723858470
transform 1 0 3083 0 -1 3605
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_1
timestamp 1723858470
transform 1 0 3083 0 1 1977
box -66 -43 450 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1723858470
transform 1 0 299 0 1 1977
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1723858470
transform 1 0 299 0 -1 3605
box -66 -43 258 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1723858470
transform 1 0 2603 0 1 1977
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_1
timestamp 1723858470
transform 1 0 2603 0 -1 3605
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1723858470
transform 1 0 491 0 1 1977
box -66 -43 2178 1671
<< labels >>
flabel metal2 0 1162 156 1308 0 FreeSans 800 0 0 0 avdd
port 4 nsew
flabel metal1 1 2530 263 2638 0 FreeSans 800 0 0 0 dvdd
port 6 nsew
flabel metal1 0 3479 263 3627 0 FreeSans 800 0 0 0 dvss
port 7 nsew
flabel metal1 2 2041 182 2130 0 FreeSans 800 0 0 0 on
port 8 nsew
flabel metal2 0 -340 156 -194 0 FreeSans 800 0 0 0 avss
port 5 nsew
flabel metal2 3308 772 3494 972 0 FreeSans 800 0 0 0 in
port 2 nsew
flabel metal2 3308 -19 3494 180 0 FreeSans 800 0 0 0 out
port 3 nsew
<< end >>
