magic
tech sky130A
magscale 1 2
timestamp 1722433690
<< dnwell >>
rect 1187 127 3988 1461
<< nwell >>
rect 1077 1190 4097 1570
rect 1077 410 1660 1190
rect 3766 410 4097 1190
rect 1077 24 4097 410
<< mvnsubdiff >>
rect 1144 1484 4031 1504
rect 1144 1450 1224 1484
rect 3951 1450 4031 1484
rect 1144 1430 4031 1450
rect 1144 1424 1218 1430
rect 1144 170 1164 1424
rect 1198 170 1218 1424
rect 1144 164 1218 170
rect 3957 1424 4031 1430
rect 3957 170 3977 1424
rect 4011 170 4031 1424
rect 3957 164 4031 170
rect 1144 144 4031 164
rect 1144 110 1224 144
rect 3951 110 4031 144
rect 1144 90 4031 110
<< mvnsubdiffcont >>
rect 1224 1450 3951 1484
rect 1164 170 1198 1424
rect 3977 170 4011 1424
rect 1224 110 3951 144
<< locali >>
rect 1164 1450 1224 1484
rect 3951 1450 4011 1484
rect 1164 1424 4011 1450
rect 1198 1348 3977 1424
rect 1198 1263 1385 1348
rect 3826 1263 3977 1348
rect 1198 1255 3977 1263
rect 1198 1220 1566 1255
rect 3936 1220 3977 1255
rect 1198 1169 3977 1220
rect 1198 244 1385 1169
rect 1657 1098 3724 1121
rect 1657 1086 3649 1098
rect 1657 509 1693 1086
rect 1749 1036 3649 1086
rect 1749 567 1800 1036
rect 3620 567 3649 1036
rect 1749 513 3649 567
rect 3696 513 3724 1098
rect 1749 509 3724 513
rect 1657 405 3724 509
rect 1657 354 1690 405
rect 3705 354 3724 405
rect 1657 341 3724 354
rect 3826 244 3977 1169
rect 1198 170 3977 244
rect 1164 144 4011 170
rect 1164 110 1224 144
rect 3951 110 4011 144
<< viali >>
rect 1566 1220 3936 1255
rect 1693 509 1749 1086
rect 3649 513 3696 1098
rect 1690 354 3705 405
<< metal1 >>
rect 1350 1255 4017 1332
rect 1350 1220 1566 1255
rect 3936 1220 4017 1255
rect 1350 1186 4017 1220
rect 1665 1086 1772 1126
rect 1665 509 1693 1086
rect 1749 509 1772 1086
rect 2614 1074 3208 1114
rect 3324 1075 3421 1111
rect 1864 781 1913 851
rect 1665 430 1772 509
rect 1997 497 2031 930
rect 2614 905 2642 1074
rect 2774 906 2802 1074
rect 2113 781 2162 851
rect 2481 781 2530 851
rect 2889 781 2938 851
rect 2614 567 2642 698
rect 2774 567 2802 699
rect 3091 567 3127 1074
rect 3384 929 3421 1075
rect 3627 1098 3715 1116
rect 2614 533 3127 567
rect 3390 497 3418 674
rect 1997 465 3418 497
rect 3627 513 3649 1098
rect 3696 513 3715 1098
rect 3627 430 3715 513
rect 1350 405 4022 430
rect 1350 354 1690 405
rect 3705 354 4022 405
rect 1350 284 4022 354
<< metal2 >>
rect 3208 1074 3248 1566
rect 3288 1075 3324 1567
rect 1854 824 3798 923
rect 3622 676 3798 677
rect 1854 587 3798 676
use iso_switch_via  iso_switch_via_0
timestamp 1722433690
transform 1 0 1829 0 -1 -2121
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_1
timestamp 1722433690
transform 0 -1 584 -1 0 1514
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_2
timestamp 1722433690
transform 0 -1 322 -1 0 1793
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_3
timestamp 1722433690
transform 0 -1 569 -1 0 1797
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_4
timestamp 1722433690
transform 1 0 1438 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_9
timestamp 1722433690
transform 1 0 2214 0 -1 -2122
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_10
timestamp 1722433690
transform 0 -1 -105 -1 0 1509
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_11
timestamp 1722433690
transform 1 0 1212 0 -1 -2129
box 652 -2914 724 -2722
use sky130_fd_pr__nfet_g5v0d10v5_SF7DK5  XM1 paramcells
timestamp 1722433690
transform 1 0 3404 0 1 801
box -308 -347 308 347
use sky130_fd_pr__nfet_g5v0d10v5_SF7DK5  XM2
timestamp 1722433690
transform 1 0 2014 0 1 801
box -308 -347 308 347
use sky130_fd_pr__nfet_g5v0d10v5_VDJU7P  XM3 paramcells
timestamp 1722433690
transform 1 0 2709 0 1 801
box -387 -347 387 347
<< labels >>
flabel metal2 3622 587 3790 677 0 FreeSans 256 180 0 0 out
port 3 nsew
flabel metal1 1350 1186 1549 1264 0 FreeSans 480 0 0 0 vdd
port 5 nsew
flabel metal2 3623 824 3789 923 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal2 3288 1386 3324 1567 0 FreeSans 256 270 0 0 off
port 1 nsew
flabel metal2 3208 1390 3248 1566 0 FreeSans 256 270 0 0 on
port 0 nsew
flabel metal1 1350 354 1551 430 0 FreeSans 480 0 0 0 vss
port 6 nsew
<< end >>
