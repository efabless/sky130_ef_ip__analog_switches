magic
tech sky130A
magscale 1 2
timestamp 1719092366
<< pwell >>
rect -515 -758 515 758
<< mvnmos >>
rect -287 -500 -187 500
rect -129 -500 -29 500
rect 29 -500 129 500
rect 187 -500 287 500
<< mvndiff >>
rect -345 488 -287 500
rect -345 -488 -333 488
rect -299 -488 -287 488
rect -345 -500 -287 -488
rect -187 488 -129 500
rect -187 -488 -175 488
rect -141 -488 -129 488
rect -187 -500 -129 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 129 488 187 500
rect 129 -488 141 488
rect 175 -488 187 488
rect 129 -500 187 -488
rect 287 488 345 500
rect 287 -488 299 488
rect 333 -488 345 488
rect 287 -500 345 -488
<< mvndiffc >>
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
<< mvpsubdiff >>
rect -479 710 479 722
rect -479 676 -371 710
rect 371 676 479 710
rect -479 664 479 676
rect -479 614 -421 664
rect -479 -614 -467 614
rect -433 -614 -421 614
rect 421 614 479 664
rect -479 -664 -421 -614
rect 421 -614 433 614
rect 467 -614 479 614
rect 421 -664 479 -614
rect -479 -676 479 -664
rect -479 -710 -371 -676
rect 371 -710 479 -676
rect -479 -722 479 -710
<< mvpsubdiffcont >>
rect -371 676 371 710
rect -467 -614 -433 614
rect 433 -614 467 614
rect -371 -710 371 -676
<< poly >>
rect -287 572 -187 588
rect -287 538 -271 572
rect -203 538 -187 572
rect -287 500 -187 538
rect -129 572 -29 588
rect -129 538 -113 572
rect -45 538 -29 572
rect -129 500 -29 538
rect 29 572 129 588
rect 29 538 45 572
rect 113 538 129 572
rect 29 500 129 538
rect 187 572 287 588
rect 187 538 203 572
rect 271 538 287 572
rect 187 500 287 538
rect -287 -538 -187 -500
rect -287 -572 -271 -538
rect -203 -572 -187 -538
rect -287 -588 -187 -572
rect -129 -538 -29 -500
rect -129 -572 -113 -538
rect -45 -572 -29 -538
rect -129 -588 -29 -572
rect 29 -538 129 -500
rect 29 -572 45 -538
rect 113 -572 129 -538
rect 29 -588 129 -572
rect 187 -538 287 -500
rect 187 -572 203 -538
rect 271 -572 287 -538
rect 187 -588 287 -572
<< polycont >>
rect -271 538 -203 572
rect -113 538 -45 572
rect 45 538 113 572
rect 203 538 271 572
rect -271 -572 -203 -538
rect -113 -572 -45 -538
rect 45 -572 113 -538
rect 203 -572 271 -538
<< locali >>
rect -467 676 -371 710
rect 371 676 467 710
rect -467 614 -433 676
rect 433 614 467 676
rect -287 538 -271 572
rect -203 538 -187 572
rect -129 538 -113 572
rect -45 538 -29 572
rect 29 538 45 572
rect 113 538 129 572
rect 187 538 203 572
rect 271 538 287 572
rect -333 488 -299 504
rect -333 -504 -299 -488
rect -175 488 -141 504
rect -175 -504 -141 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 141 488 175 504
rect 141 -504 175 -488
rect 299 488 333 504
rect 299 -504 333 -488
rect -287 -572 -271 -538
rect -203 -572 -187 -538
rect -129 -572 -113 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 113 -572 129 -538
rect 187 -572 203 -538
rect 271 -572 287 -538
rect -467 -676 -433 -614
rect 433 -676 467 -614
rect -467 -710 -371 -676
rect 371 -710 467 -676
<< viali >>
rect -271 538 -203 572
rect -113 538 -45 572
rect 45 538 113 572
rect 203 538 271 572
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect -271 -572 -203 -538
rect -113 -572 -45 -538
rect 45 -572 113 -538
rect 203 -572 271 -538
<< metal1 >>
rect -283 572 -191 578
rect -283 538 -271 572
rect -203 538 -191 572
rect -283 532 -191 538
rect -125 572 -33 578
rect -125 538 -113 572
rect -45 538 -33 572
rect -125 532 -33 538
rect 33 572 125 578
rect 33 538 45 572
rect 113 538 125 572
rect 33 532 125 538
rect 191 572 283 578
rect 191 538 203 572
rect 271 538 283 572
rect 191 532 283 538
rect -339 488 -293 500
rect -339 -488 -333 488
rect -299 -488 -293 488
rect -339 -500 -293 -488
rect -181 488 -135 500
rect -181 -488 -175 488
rect -141 -488 -135 488
rect -181 -500 -135 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 135 488 181 500
rect 135 -488 141 488
rect 175 -488 181 488
rect 135 -500 181 -488
rect 293 488 339 500
rect 293 -488 299 488
rect 333 -488 339 488
rect 293 -500 339 -488
rect -283 -538 -191 -532
rect -283 -572 -271 -538
rect -203 -572 -191 -538
rect -283 -578 -191 -572
rect -125 -538 -33 -532
rect -125 -572 -113 -538
rect -45 -572 -33 -538
rect -125 -578 -33 -572
rect 33 -538 125 -532
rect 33 -572 45 -538
rect 113 -572 125 -538
rect 33 -578 125 -572
rect 191 -538 283 -532
rect 191 -572 203 -538
rect 271 -572 283 -538
rect 191 -578 283 -572
<< properties >>
string FIXED_BBOX -450 -693 450 693
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5.0 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
