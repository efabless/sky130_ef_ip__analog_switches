magic
tech sky130A
magscale 1 2
timestamp 1722434346
<< psubdiff >>
rect 491 1640 515 1724
rect 3454 1640 3478 1724
<< psubdiffcont >>
rect 515 1640 3454 1724
<< locali >>
rect 2566 3229 2629 3295
rect 2879 3275 3095 3283
rect 2879 3230 2890 3275
rect 3085 3230 3095 3275
rect 2879 3221 3095 3230
rect 756 2379 996 2392
rect 756 2337 770 2379
rect 982 2337 996 2379
rect 756 2324 996 2337
rect 2444 2347 2684 2353
rect 2444 2295 2460 2347
rect 2668 2295 2684 2347
rect 2444 2287 2684 2295
rect 2851 2348 3058 2354
rect 2851 2296 2867 2348
rect 2851 2288 3058 2296
rect 402 2048 458 2056
rect 402 1964 410 2048
rect 448 1994 458 2048
rect 448 1964 492 1994
rect 402 1960 492 1964
rect 402 1954 458 1960
rect 499 1640 515 1724
rect 3454 1640 3470 1724
<< viali >>
rect 2890 3230 3085 3275
rect 770 2337 982 2379
rect 3157 2363 3207 2499
rect 2460 2295 2668 2347
rect 2867 2296 3058 2348
rect 410 1964 448 2048
rect 1009 1640 1199 1724
<< metal1 >>
rect 350 3604 651 3627
rect 350 3559 3461 3604
rect 350 3538 1011 3559
rect 350 3479 651 3538
rect 1001 3430 1011 3538
rect 1198 3538 3461 3559
rect 1198 3430 1208 3538
rect 1001 3420 1208 3430
rect 2869 3275 3111 3283
rect 2869 3230 2890 3275
rect 3085 3230 3111 3275
rect 2869 3221 3111 3230
rect 615 2903 837 2916
rect 615 2868 627 2903
rect 491 2730 627 2868
rect 615 2677 627 2730
rect 826 2868 837 2903
rect 1804 2903 2027 2916
rect 1804 2868 1816 2903
rect 826 2730 1816 2868
rect 826 2677 837 2730
rect 615 2666 837 2677
rect 1804 2678 1816 2730
rect 2013 2868 2027 2903
rect 2013 2730 3464 2868
rect 2013 2678 2027 2730
rect 1804 2666 2027 2678
rect 351 2581 651 2638
rect 351 2530 613 2581
rect 1395 2499 3214 2515
rect 1395 2479 3157 2499
rect 756 2379 996 2392
rect 352 2365 639 2366
rect 756 2365 770 2379
rect 352 2337 770 2365
rect 982 2365 996 2379
rect 1395 2365 1431 2479
rect 982 2337 1431 2365
rect 3150 2363 3157 2479
rect 3207 2363 3214 2499
rect 352 2329 1431 2337
rect 2444 2347 2684 2353
rect 352 2277 639 2329
rect 756 2324 996 2329
rect 2444 2295 2460 2347
rect 2668 2295 2684 2347
rect 2444 2287 2684 2295
rect 2851 2348 3058 2354
rect 2851 2296 2867 2348
rect 3150 2345 3214 2363
rect 2851 2288 3058 2296
rect 398 2048 3468 2056
rect 398 1964 410 2048
rect 448 1980 3468 2048
rect 448 1964 496 1980
rect 398 1954 496 1964
rect 996 1724 1213 1735
rect 996 1640 1009 1724
rect 1199 1640 1213 1724
rect 996 1630 1213 1640
rect 350 1302 837 1308
rect 350 1169 624 1302
rect 830 1169 837 1302
rect 350 1162 837 1169
rect 1805 1301 2027 1308
rect 1805 1170 1814 1301
rect 2019 1170 2027 1301
rect 1805 1162 2027 1170
rect 350 260 773 406
<< via1 >>
rect 1011 3430 1198 3559
rect 627 2677 826 2903
rect 1816 2678 2013 2903
rect 1009 1640 1199 1724
rect 624 1169 830 1302
rect 1814 1170 2019 1301
<< metal2 >>
rect 1001 3559 1208 3568
rect 1001 3430 1011 3559
rect 1198 3430 1208 3559
rect 615 2903 837 2916
rect 615 2677 627 2903
rect 826 2677 837 2903
rect 615 1302 837 2677
rect 1001 1724 1208 3430
rect 1804 2903 2027 2916
rect 1804 2678 1816 2903
rect 2013 2678 2027 2903
rect 1804 2666 2027 2678
rect 1001 1640 1009 1724
rect 1199 1640 1208 1724
rect 1001 1630 1208 1640
rect 615 1169 624 1302
rect 830 1169 837 1302
rect 615 1162 837 1169
rect 1805 1301 2027 2666
rect 2883 2471 2931 3252
rect 2626 2423 3181 2471
rect 2418 2282 2468 2353
rect 2626 2283 2674 2423
rect 2801 2287 2883 2359
rect 2958 2287 3006 2295
rect 2801 2232 2851 2287
rect 2631 2182 2851 2232
rect 2631 1540 2671 2182
rect 3133 2130 3181 2423
rect 2711 2082 3181 2130
rect 2711 1543 2747 2082
rect 1805 1170 1814 1301
rect 2019 1170 2027 1301
rect 1805 1162 2027 1170
rect 3218 800 3516 899
rect 3219 563 3516 653
use iso_switch_via  iso_switch_via_0
timestamp 1722433690
transform 0 1 5797 1 0 2564
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_1
timestamp 1722433690
transform 0 1 5380 1 0 1630
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_2
timestamp 1722433690
transform 0 1 5797 1 0 1635
box 652 -2914 724 -2722
use minimum_analog_switch  minimum_analog_switch_0
timestamp 1722433690
transform 1 0 -577 0 1 -24
box 1077 24 4097 1570
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1722433690
transform 1 0 3083 0 -1 3605
box -66 -43 450 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1722433690
transform 1 0 3083 0 1 1977
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1722433690
transform 1 0 3275 0 1 1977
box -66 -43 258 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1722433690
transform 1 0 2603 0 1 1977
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_1
timestamp 1722433690
transform 1 0 2603 0 -1 3605
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1722433690
transform 1 0 491 0 1 1977
box -66 -43 2178 1671
<< labels >>
flabel metal1 351 2530 613 2638 0 FreeSans 800 0 0 0 dvdd
port 6 nsew
flabel metal1 350 3479 613 3627 0 FreeSans 800 0 0 0 dvss
port 7 nsew
flabel metal1 352 2277 532 2366 0 FreeSans 800 0 0 0 on
port 8 nsew
flabel metal2 3330 800 3516 899 0 FreeSans 800 0 0 0 in
port 2 nsew
flabel metal1 350 260 506 406 0 FreeSans 800 0 0 0 avss
port 5 nsew
flabel metal1 350 1162 506 1308 0 FreeSans 800 0 0 0 avdd
port 4 nsew
flabel metal2 3330 563 3516 653 0 FreeSans 800 0 0 0 out
port 3 nsew
<< end >>
