magic
tech sky130A
timestamp 1719092895
<< metal1 >>
rect 306 -1245 382 -1241
rect 306 -1453 310 -1245
rect 377 -1453 382 -1245
rect 306 -1457 382 -1453
<< via1 >>
rect 310 -1453 377 -1245
<< metal2 >>
rect 306 -1245 382 -1241
rect 306 -1453 310 -1245
rect 377 -1453 382 -1245
rect 306 -1457 382 -1453
<< end >>
