magic
tech sky130A
magscale 1 2
timestamp 1722433690
<< pwell >>
rect -387 -347 387 347
<< mvnmos >>
rect -129 -50 -29 50
rect 29 -50 129 50
<< mvndiff >>
rect -187 38 -129 50
rect -187 -38 -175 38
rect -141 -38 -129 38
rect -187 -50 -129 -38
rect -29 38 29 50
rect -29 -38 -17 38
rect 17 -38 29 38
rect -29 -50 29 -38
rect 129 38 187 50
rect 129 -38 141 38
rect 175 -38 187 38
rect 129 -50 187 -38
<< mvndiffc >>
rect -175 -38 -141 38
rect -17 -38 17 38
rect 141 -38 175 38
<< mvpsubdiff >>
rect -321 269 321 281
rect -321 235 -213 269
rect 213 235 321 269
rect -321 223 321 235
rect -321 173 -263 223
rect -321 -173 -309 173
rect -275 -173 -263 173
rect 263 173 321 223
rect -321 -223 -263 -173
rect 263 -173 275 173
rect 309 -173 321 173
rect 263 -223 321 -173
rect -321 -235 321 -223
rect -321 -269 -213 -235
rect 213 -269 321 -235
rect -321 -281 321 -269
<< mvpsubdiffcont >>
rect -213 235 213 269
rect -309 -173 -275 173
rect 275 -173 309 173
rect -213 -269 213 -235
<< poly >>
rect -129 131 -29 147
rect -129 97 -113 131
rect -45 97 -29 131
rect -129 50 -29 97
rect 29 131 129 147
rect 29 97 45 131
rect 113 97 129 131
rect 29 50 129 97
rect -129 -97 -29 -50
rect -129 -131 -113 -97
rect -45 -131 -29 -97
rect -129 -147 -29 -131
rect 29 -97 129 -50
rect 29 -131 45 -97
rect 113 -131 129 -97
rect 29 -147 129 -131
<< polycont >>
rect -113 97 -45 131
rect 45 97 113 131
rect -113 -131 -45 -97
rect 45 -131 113 -97
<< locali >>
rect -309 235 -213 269
rect 213 235 309 269
rect -309 173 -275 235
rect 275 173 309 235
rect -129 97 -113 131
rect -45 97 -29 131
rect 29 97 45 131
rect 113 97 129 131
rect -175 38 -141 54
rect -175 -54 -141 -38
rect -17 38 17 54
rect -17 -54 17 -38
rect 141 38 175 54
rect 141 -54 175 -38
rect -129 -131 -113 -97
rect -45 -131 -29 -97
rect 29 -131 45 -97
rect 113 -131 129 -97
rect -309 -235 -275 -173
rect 275 -235 309 -173
rect -309 -269 -213 -235
rect 213 -269 309 -235
<< viali >>
rect -113 97 -45 131
rect 45 97 113 131
rect -175 -38 -141 38
rect -17 -38 17 38
rect 141 -38 175 38
rect -113 -131 -45 -97
rect 45 -131 113 -97
<< metal1 >>
rect -125 131 -33 137
rect -125 97 -113 131
rect -45 97 -33 131
rect -125 91 -33 97
rect 33 131 125 137
rect 33 97 45 131
rect 113 97 125 131
rect 33 91 125 97
rect -181 38 -135 50
rect -181 -38 -175 38
rect -141 -38 -135 38
rect -181 -50 -135 -38
rect -23 38 23 50
rect -23 -38 -17 38
rect 17 -38 23 38
rect -23 -50 23 -38
rect 135 38 181 50
rect 135 -38 141 38
rect 175 -38 181 38
rect 135 -50 181 -38
rect -125 -97 -33 -91
rect -125 -131 -113 -97
rect -45 -131 -33 -97
rect -125 -137 -33 -131
rect 33 -97 125 -91
rect 33 -131 45 -97
rect 113 -131 125 -97
rect 33 -137 125 -131
<< properties >>
string FIXED_BBOX -292 -252 292 252
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.5 l 0.5 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8  sky130_fd_pr__nfet_01v8_lvt sky130_fd_pr__nfet_01v8_hvt  sky130_fd_pr__nfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
