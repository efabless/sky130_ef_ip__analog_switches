** sch_path: /home/tim/gits/sky130_ef_ip__analog_switches/xschem/isolated_switch_large.sch
.subckt isolated_switch_large avss on out in avdd dvdd dvss off
*.PININFO on:I avss:B out:B in:B avdd:B dvdd:B dvss:B off:I
x2 on dvdd dvss dvss avdd avdd net1 sky130_fd_sc_hvl__lsbuflv2hv_1
XD1 dvss on sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
x1 net1 net2 avss out in avdd net3 isolated_switch_3
x3 off dvdd dvss dvss avdd avdd net3 sky130_fd_sc_hvl__lsbuflv2hv_1
XD2 dvss off sky130_fd_pr__diode_pw2nd_05v5 area=2.025e11 perim=1.8e6
x4 net1 dvss dvss avdd avdd net2 sky130_fd_sc_hvl__inv_1
.ends

* expanding   symbol:  isolated_switch_3.sym # of pins=7
** sym_path: /home/tim/gits/sky130_ef_ip__analog_switches/xschem/isolated_switch_3.sym
** sch_path: /home/tim/gits/sky130_ef_ip__analog_switches/xschem/isolated_switch_3.sch
.subckt isolated_switch_3 on off vss out in vdd shunt
*.PININFO on:I out:B vdd:B vss:B in:B off:I shunt:I
XM1 in on net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=12 nf=6 m=1
XM2 in off net1 vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=24 nf=12 m=1
XM11 net1 on out vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=12 nf=6 m=1
XM12 net1 off out vdd sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=24 nf=12 m=1
XM17 vss shunt net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends

.end
