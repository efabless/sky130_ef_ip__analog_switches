magic
tech sky130A
magscale 1 2
timestamp 1716596057
<< dnwell >>
rect 687 -653 5284 1461
rect 687 -659 2073 -653
<< nwell >>
rect 577 1255 5393 1570
rect 577 -447 773 1255
rect 5078 -447 5393 1255
rect 577 -762 5393 -447
<< mvnsubdiff >>
rect 644 1484 5327 1504
rect 644 1450 724 1484
rect 5247 1450 5327 1484
rect 644 1430 5327 1450
rect 644 1424 718 1430
rect 644 -616 664 1424
rect 698 -616 718 1424
rect 644 -622 718 -616
rect 5253 1424 5327 1430
rect 5253 -616 5273 1424
rect 5307 -616 5327 1424
rect 5253 -622 5327 -616
rect 644 -642 5327 -622
rect 644 -676 724 -642
rect 5247 -676 5327 -642
rect 644 -696 5327 -676
<< mvnsubdiffcont >>
rect 724 1450 5247 1484
rect 664 -616 698 1424
rect 5273 -616 5307 1424
rect 724 -676 5247 -642
<< locali >>
rect 664 1450 724 1484
rect 5247 1450 5307 1484
rect 664 1424 5307 1450
rect 698 1348 5273 1424
rect 698 1263 885 1348
rect 3560 1276 5028 1286
rect 698 1255 2954 1263
rect 698 1220 1066 1255
rect 2929 1220 2954 1255
rect 698 1169 2954 1220
rect 3560 1230 3582 1276
rect 5010 1230 5028 1276
rect 3560 1196 5028 1230
rect 698 -542 885 1169
rect 3560 -407 5063 -345
rect 3560 -444 3603 -407
rect 4840 -444 5063 -407
rect 3560 -462 5063 -444
rect 5122 -542 5273 1348
rect 698 -616 5273 -542
rect 664 -642 5307 -616
rect 664 -676 724 -642
rect 5247 -676 5307 -642
<< viali >>
rect 1066 1220 2929 1255
rect 3582 1230 5010 1276
rect 3603 -444 4840 -407
<< metal1 >>
rect 3194 1390 3261 1566
rect 850 1264 3152 1332
rect 849 1255 3152 1264
rect 849 1220 1066 1255
rect 2929 1220 3152 1255
rect 849 1186 3152 1220
rect 1035 1046 1285 1092
rect 1619 1046 2185 1095
rect 2519 1046 2769 1095
rect 3208 1074 3248 1390
rect 3334 1386 3402 1567
rect 1065 564 1093 1046
rect 1224 564 1252 1046
rect 1649 567 1677 1046
rect 1807 567 1835 1046
rect 1967 567 1995 1046
rect 2125 567 2153 1046
rect 2549 567 2577 1046
rect 2709 567 2737 1046
rect 3348 574 3384 1386
rect 3458 1276 5081 1332
rect 3458 1230 3582 1276
rect 5010 1230 5081 1276
rect 3458 1186 5081 1230
rect 1035 518 1285 564
rect 1619 518 2185 567
rect 2519 518 2769 567
rect 1065 291 1093 518
rect 1224 291 1252 518
rect 1649 291 1677 518
rect 1807 291 1835 518
rect 1967 291 1995 518
rect 2125 291 2153 518
rect 2549 291 2577 518
rect 2709 291 2737 518
rect 3139 512 3247 517
rect 3139 501 3322 512
rect 3139 327 3148 501
rect 3238 327 3322 501
rect 3139 312 3322 327
rect 1035 245 1285 291
rect 1619 245 1677 291
rect 1679 245 1835 291
rect 1837 245 1995 291
rect 1996 245 2185 291
rect 2519 245 2577 291
rect 2580 245 2737 291
rect 2738 245 2769 291
rect 1065 -237 1093 245
rect 1224 -237 1252 245
rect 1649 -235 1677 245
rect 1807 -235 1835 245
rect 1967 -235 1995 245
rect 2125 -235 2153 245
rect 1035 -283 1285 -237
rect 1619 -283 2185 -235
rect 2549 -237 2577 245
rect 2709 -237 2737 245
rect 2519 -283 2577 -237
rect 2580 -283 2737 -237
rect 2738 -283 2769 -237
rect 2549 -284 2577 -283
rect 3139 -356 3247 312
rect 3352 238 3380 574
rect 3344 -260 3386 238
rect 3778 -251 3806 1067
rect 4170 1029 4420 1075
rect 4204 568 4232 1029
rect 4362 568 4390 1029
rect 4170 519 4420 568
rect 4204 289 4232 519
rect 4362 289 4390 519
rect 4170 243 4203 289
rect 4204 243 4359 289
rect 4362 243 4420 289
rect 4204 -221 4232 243
rect 4362 -221 4390 243
rect 3352 -284 3380 -260
rect 4170 -267 4203 -221
rect 4204 -267 4359 -221
rect 4362 -267 4420 -221
rect 4788 -251 4816 1067
rect 832 -407 5063 -356
rect 832 -444 3603 -407
rect 4840 -444 5063 -407
rect 832 -502 5063 -444
<< via1 >>
rect 3148 327 3238 501
<< metal2 >>
rect 964 1074 4869 1114
rect 4886 1016 5062 1023
rect 965 824 5062 1016
rect 4886 823 5062 824
rect 965 584 4924 776
rect 3139 501 3320 509
rect 3139 327 3148 501
rect 3238 327 3320 501
rect 3139 319 3320 327
rect 3410 235 3607 584
rect 965 43 4832 235
rect 4886 -17 5062 -9
rect 965 -209 5062 -17
rect 964 -305 4864 -265
use iso_switch_via  iso_switch_via_0
timestamp 1716573125
transform 0 -1 -917 -1 0 397
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_1
timestamp 1716573125
transform 1 0 1373 0 -1 -1900
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_2
timestamp 1716573125
transform -1 0 4986 0 -1 -1914
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_3
timestamp 1716573125
transform 1 0 1533 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_4
timestamp 1716573125
transform 1 0 1211 0 -1 -2124
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_5
timestamp 1716573125
transform 1 0 897 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_6
timestamp 1716573125
transform 1 0 633 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_7
timestamp 1716573125
transform 1 0 471 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_8
timestamp 1716573125
transform 1 0 1797 0 -1 -1904
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_9
timestamp 1716573125
transform 1 0 2113 0 -1 -1904
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_10
timestamp 1716573125
transform 1 0 1955 0 -1 -1904
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_11
timestamp 1716573125
transform 1 0 1053 0 -1 -1898
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_12
timestamp 1716573125
transform 1 0 1053 0 1 2925
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_13
timestamp 1716573125
transform 1 0 1371 0 1 2925
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_14
timestamp 1716573125
transform 1 0 1211 0 1 2715
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_15
timestamp 1716573125
transform 1 0 1529 0 1 2715
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_16
timestamp 1716573125
transform 1 0 1795 0 1 2933
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_17
timestamp 1716573125
transform 1 0 313 0 1 2705
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_18
timestamp 1716573125
transform 1 0 1953 0 1 2931
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_19
timestamp 1716573125
transform 1 0 2113 0 1 2935
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_20
timestamp 1716573125
transform 1 0 629 0 1 2709
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_21
timestamp 1716573125
transform 1 0 469 0 1 2709
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_22
timestamp 1716573125
transform 1 0 895 0 1 2709
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_23
timestamp 1716573125
transform -1 0 5146 0 -1 -2120
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_24
timestamp 1716573125
transform -1 0 4824 0 -1 -2120
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_25
timestamp 1716573125
transform -1 0 5410 0 -1 -2124
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_26
timestamp 1716573125
transform -1 0 4560 0 -1 -1916
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_27
timestamp 1716573125
transform -1 0 4402 0 -1 -1914
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_28
timestamp 1716573125
transform -1 0 5146 0 1 2723
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_29
timestamp 1716573125
transform -1 0 5570 0 -1 -2124
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_30
timestamp 1716573125
transform -1 0 5568 0 1 2721
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_31
timestamp 1716573125
transform -1 0 5412 0 1 2723
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_32
timestamp 1716573125
transform -1 0 4828 0 1 2721
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_33
timestamp 1716573125
transform -1 0 4984 0 1 2937
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_34
timestamp 1716573125
transform -1 0 4402 0 1 2935
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_35
timestamp 1716573125
transform -1 0 4562 0 1 2935
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_36
timestamp 1716573125
transform -1 0 3974 0 1 3234
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_37
timestamp 1716573125
transform -1 0 4134 0 1 3235
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_38
timestamp 1716573125
transform 1 0 313 0 -1 -2126
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_40
timestamp 1716573125
transform 0 -1 971 -1 0 397
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_41
timestamp 1716573125
transform 0 -1 -1671 -1 0 1799
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_42
timestamp 1716573125
transform 0 -1 1979 -1 0 399
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_43
timestamp 1716573125
transform 0 1 5976 1 0 410
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_44
timestamp 1716573125
transform 0 -1 1487 -1 0 1799
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_45
timestamp 1716573125
transform 0 -1 -151 -1 0 1799
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_47
timestamp 1716573125
transform 0 -1 -163 -1 0 987
box 652 -2914 724 -2722
use iso_switch_via  iso_switch_via_53
timestamp 1716573125
transform 0 -1 571 -1 0 397
box 652 -2914 724 -2722
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  sky130_fd_pr__nfet_g5v0d10v5_EJGQJV_0 paramcells
timestamp 1716587504
transform -1 0 3366 0 1 412
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_E7BQJJ  XM1 paramcells
timestamp 1716587504
transform -1 0 4295 0 1 797
box -357 -458 357 458
use sky130_fd_pr__pfet_g5v0d10v5_KLHCT5  XM2 paramcells
timestamp 1716587504
transform 1 0 1902 0 1 4
box -545 -497 545 497
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM3 paramcells
timestamp 1716587504
transform -1 0 4800 0 1 797
box -278 -458 278 458
use sky130_fd_pr__pfet_g5v0d10v5_KL97Y6  XM4 paramcells
timestamp 1716587504
transform 1 0 1160 0 1 4
box -387 -497 387 497
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM5
timestamp 1716587504
transform -1 0 3790 0 1 797
box -278 -458 278 458
use sky130_fd_pr__pfet_g5v0d10v5_KL97Y6  XM6
timestamp 1716587504
transform 1 0 2644 0 1 4
box -387 -497 387 497
use sky130_fd_pr__nfet_g5v0d10v5_E7BQJJ  XM11
timestamp 1716587504
transform -1 0 4295 0 1 11
box -357 -458 357 458
use sky130_fd_pr__pfet_g5v0d10v5_KLHCT5  XM12
timestamp 1716587504
transform 1 0 1902 0 1 808
box -545 -497 545 497
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM13
timestamp 1716587504
transform -1 0 4800 0 1 11
box -278 -458 278 458
use sky130_fd_pr__pfet_g5v0d10v5_KL97Y6  XM14
timestamp 1716587504
transform 1 0 1160 0 1 808
box -387 -497 387 497
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM15
timestamp 1716587504
transform -1 0 3790 0 1 11
box -278 -458 278 458
use sky130_fd_pr__pfet_g5v0d10v5_KL97Y6  XM16
timestamp 1716587504
transform 1 0 2644 0 1 808
box -387 -497 387 497
<< labels >>
flabel metal2 4886 -209 5062 -9 0 FreeSans 256 180 0 0 out
port 3 nsew
flabel metal1 849 1186 1049 1264 0 FreeSans 256 0 0 0 vdd
port 5 nsew
flabel metal2 4886 823 5062 1023 0 FreeSans 256 0 0 0 in
port 4 nsew
flabel metal1 832 -463 1032 -356 0 FreeSans 256 180 0 0 vss
port 2 nsew
flabel metal1 3194 1390 3261 1566 0 FreeSans 256 270 0 0 on
port 0 nsew
flabel metal1 3334 1386 3402 1567 0 FreeSans 256 270 0 0 off
port 1 nsew
<< end >>
